`timescale 1ns / 1ps

module keccak_f1600_tb;

    // DUT signals
    reg          clk;
    reg          rst_n;
    reg          start;
    reg  [1599:0] state_in;
    wire [1599:0] state_out;
    wire         ready;
    wire         done;

    // Instantiate DUT
    keccak_f1600 uut (
        .clk       (clk),
        .rst_n     (rst_n),
        .start     (start),
        .state_in  (state_in),
        .state_out (state_out),
        .ready     (ready),
        .done      (done)
    );

    // 10 ns clock period
    always #5 clk = ~clk;

    // Reference vectors: 2 test cases x 25 lanes = 50 entries
    // Generated by gen_f1600_vectors.cpp
    reg [63:0] expected_lanes [0:49];

    integer i, errors;
    reg [1599:0] expected_state;

    // Display all 25 lanes
    task display_state;
        input [1599:0] s;
        integer k;
        begin
            for (k = 0; k < 25; k = k + 1)
                $display("  Lane[%2d] = %h", k, s[k*64 +: 64]);
        end
    endtask

    // Build 1600-bit expected state from lane array starting at base index
    task build_expected;
        input integer base;
        integer k;
        begin
            expected_state = 1600'd0;
            for (k = 0; k < 25; k = k + 1)
                expected_state[k*64 +: 64] = expected_lanes[base + k];
        end
    endtask

    // Compare state_out with expected and report
    task check_output;
        input integer test_num;
        input integer base;
        reg pass;
        integer k;
        begin
            build_expected(base);
            pass = 1;

            if (state_out !== expected_state) begin
                $display("FAIL: Test %0d", test_num);
                for (k = 0; k < 25; k = k + 1) begin
                    if (state_out[k*64 +: 64] !== expected_lanes[base + k])
                        $display("  Lane[%2d]: expected %h, got %h",
                                 k, expected_lanes[base + k], state_out[k*64 +: 64]);
                end
                errors = errors + 1;
                pass = 0;
            end

            if (pass)
                $display("PASS: Test %0d", test_num);
        end
    endtask

    // Run one permutation: set state_in, pulse start, wait for result
    task run_permutation;
        input [1599:0] input_state;
        begin
            state_in = input_state;
            @(posedge clk);
            start <= 1;
            @(posedge clk);
            start <= 0;

            // Wait for done (registered: state_out is valid when done is high)
            wait (done == 1);
            #1;
        end
    endtask

    initial begin
        $dumpfile("keccak_f1600_tb.vcd");
        $dumpvars(0, keccak_f1600_tb);

        $readmemh("f1600_vectors.hex", expected_lanes);

        clk   = 0;
        rst_n = 0;
        start = 0;
        state_in = 1600'd0;
        errors = 0;

        // ============================================
        // Reset
        // ============================================
        #20;
        rst_n = 1;
        @(posedge clk);
        #1;

        if (!ready) begin
            $display("FAIL: ready should be high after reset");
            errors = errors + 1;
        end else
            $display("OK: ready is high after reset");

        // ============================================
        // Test 1: keccak_f1600(all-zeros)
        // ============================================
        $display("\n=== Test 1: All-zero state ===");
        run_permutation(1600'd0);

        // Verify ready returned high
        if (!ready) begin
            $display("FAIL: ready should be high after completion");
            errors = errors + 1;
        end

        check_output(1, 0);

        // ============================================
        // Test 2: keccak_f1600(lane0 = 0xDEADBEEFCAFEBABE)
        // ============================================
        $display("\n=== Test 2: Non-zero state ===");
        begin : test2_setup
            reg [1599:0] t2_in;
            t2_in = 1600'd0;
            t2_in[63:0] = 64'hDEADBEEFCAFEBABE;
            run_permutation(t2_in);
        end

        check_output(2, 25);

        // ============================================
        // Test 3: Back-to-back operation
        // Run all-zeros again immediately to verify
        // the module can be reused without extra delay.
        // ============================================
        $display("\n=== Test 3: Back-to-back (repeat all-zeros) ===");
        run_permutation(1600'd0);
        check_output(3, 0);

        // ============================================
        // Summary
        // ============================================
        $display("\n=== Summary ===");
        if (errors == 0)
            $display("ALL TESTS PASSED");
        else
            $display("FAILED: %0d error(s)", errors);

        $finish;
    end

endmodule
