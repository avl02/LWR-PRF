// UPDATE TO USE SHAKE-256 - CURRENTLY A TEMPLATE THAT READS PLACEHOLDER VALUES
module hash_to_vector #(
    parameter N_LWR = 445,
    parameter N = 2048,
    parameter ELEM_WIDTH = 12
) (
    input wire clk,
    input wire rst_n,
    input wire start,
    input wire [63:0] nonce,      // Not used in stub version
    input wire [63:0] index,      // Not used in stub version

    output reg [ELEM_WIDTH-1:0] hash_out,
    output reg [$clog2(N_LWR)-1:0] hash_idx,
    output reg hash_valid,
    output reg hash_last,
    output reg done
);

    // Memory to store pre-computed hash values from Python
    reg [ELEM_WIDTH-1:0] hash_mem [0:N_LWR-1];

    // Load hash vector from file (generated by Python script)
    initial begin
        $readmemh("hash_vector.mem", hash_mem);
    end

    // Counter to iterate through hash values
    reg [$clog2(N_LWR)-1:0] counter;

    // State machine
    localparam IDLE = 2'b00;
    localparam STREAMING = 2'b01;
    localparam DONE_STATE = 2'b10;

    reg [1:0] state;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            counter <= 0;
            hash_out <= 0;
            hash_idx <= 0;
            hash_valid <= 0;
            hash_last <= 0;
            done <= 0;
        end else begin
            case (state)
                IDLE: begin
                    hash_valid <= 0;
                    hash_last <= 0;
                    done <= 0;

                    if (start) begin
                        counter <= 0;
                        state <= STREAMING;
                    end
                end

                STREAMING: begin
                    // Output current hash value
                    hash_out <= hash_mem[counter];
                    hash_idx <= counter;
                    hash_valid <= 1;
                    hash_last <= (counter == N_LWR - 1);

                    if (counter == N_LWR - 1) begin
                        state <= DONE_STATE;
                        done <= 1;
                    end else begin
                        counter <= counter + 1;
                    end
                end

                DONE_STATE: begin
                    hash_valid <= 0;
                    hash_last <= 0;
                    // Stay in done state until reset or new start
                    if (start) begin
                        counter <= 0;
                        done <= 0;
                        state <= STREAMING;
                    end
                end

                default: state <= IDLE;
            endcase
        end
    end

endmodule
